localparam MOV = 6'b000000;
localparam JMP = 6'b000001;
localparam SLP = 6'b000010;
localparam HLT = 6'b000011;

localparam ADD = 6'b000100;
localparam SUB = 6'b000101;
localparam MUL = 6'b000110;
localparam DIV = 6'b000111;
localparam LSHIFT = 6'b001000;
localparam RSHIFT = 6'b001001;
localparam ROTL = 6'b001010;
localparam ROTR = 6'b001011;
localparam AND = 6'b001100;
localparam OR = 6'b001101;
localparam XOR = 6'b001110;
localparam NAND = 6'b001111;
localparam NOR = 6'b010000;
localparam XNOR = 6'b010001;
localparam GRT = 6'b010010;
localparam EQ = 6'b010011;