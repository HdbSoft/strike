//-----------------------------------
// The strike project, open source
// 4-bit processor written in
// Verilog and Cython
//
// strike.v - Main file
//-----------------------------------

module strike_CPU();

initial begin
	$display ("Hello, world!");
	$finish;
end


endmodule
