localparam MOV = 8'b00000000;
localparam JMP = 8'b00000001;
localparam SLP = 8'b00000010;

localparam ADD = 8'b00000011;
localparam SUB = 8'b00000100;
localparam MUL = 8'b00000101;
localparam DIV = 8'b00000110;
localparam LSHIFT = 8'b00000111;
localparam RSHIFT = 8'b00001000;
localparam ROTL = 8'b00001001;
localparam ROTR = 8'b00001010;
localparam AND = 8'b00001011;
localparam OR = 8'b00001100;
localparam XOR = 8'b00001101;
localparam NAND = 8'b00001110;
localparam NOR = 8'b00001111;
localparam XNOR = 8'b00010000;
localparam GRT = 8'b00010001;
localparam EQ = 8'b00010010;